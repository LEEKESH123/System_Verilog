class parent;
	rand int a;

	function void print();
	$display("a=%p",a);
	endfunction 

endclass

class child;
	rand int b;
	
endclass

module tb;
	

endmodule
